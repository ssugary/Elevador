-- ainda falta implementar :p