library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.Tipos_Elevadores.all;

entity Controlador is               -- 80% disso foi gpt, n�o confio (estava sem tempo e fiz isso para ter uma base :p )
    port (
        CLK             : in  std_logic;
        RESET           : in  std_logic;
        
        -- INs do Sistema / Supervisor
        andar_atual_in  : in  std_logic_vector(4 downto 0);      -- LIDO do sensor de andar
        andar_destino_in: in  std_logic_vector(4 downto 0);      -- ESCOLHIDO pelo Supervisor_Global/Unico
        direcao_req_in  : in  std_logic;                         -- DIRE��O ESCOLHIDA pelo Supervisor
        door_closed_in  : in  std_logic;                         -- LIDO do m�dulo 'porta.vhd'
        
        -- IN/OUT do Teclado (Para LIMPAR chamadas internas)
        botoes_pendentes_in  : in  std_logic_vector(31 downto 0); -- LIDO do 'keyboard.vhd'
        botoes_pendentes_out : out std_logic_vector(31 downto 0); -- ENVIADO de volta ao 'keyboard.vhd'
        
        -- OUTs para o Hardware (Porta e Motor)
        start_close_out : out std_logic;                         -- ENVIADO para 'porta.vhd'
        motor_enable_out: out std_logic;                         -- LIGAR/DESLIGAR motor
        move_up_out     : out std_logic;                         -- SENTIDO para motor (Subir)
        move_down_out   : out std_logic                          -- SENTIDO para motor (Descer)
    );
    end Controlador;
    architecture Behavioral of Controlador is
    -- Defini��o dos estados da FSM
    signal estado_atual, proximo_estado : t_estado;
    
    -- Sinais auxiliares para limpar o bot�o
    signal botoes_temp : std_logic_vector(31 downto 0);

begin
    
    -- ---------------------------------------
    -- Processo 1: M�quina de Estados (Registrador de Estado)
    -- ---------------------------------------
    process (CLK, RESET) is
    begin
        if RESET = '1' then
            estado_atual <= IDLE;
            botoes_temp  <= (others => '0');
        elsif rising_edge(CLK) then
            estado_atual <= proximo_estado;
            botoes_temp  <= botoes_pendentes_in;
        end if;
    end process;
    
    botoes_pendentes_out <= botoes_temp; -- Passa os pedidos para o teclado, exceto quando limpa

    -- ---------------------------------------
    -- Processo 2: L�gica Combinacional (Pr�ximo Estado e Sa�das)
    -- ---------------------------------------
    process (estado_atual, andar_atual_in, andar_destino_in, direcao_req_in, door_closed_in, botoes_pendentes_in, botoes_temp) is
        -- Convers�o para Integer, pois � mais f�cil de comparar
        variable atual_int    : integer;
        variable destino_int  : integer;
    begin
        -- Default: Nenhuma a��o
        proximo_estado   <= estado_atual;
        motor_enable_out <= '0';
        move_up_out      <= '0';
        move_down_out    <= '0';
        start_close_out  <= '0';

        atual_int   := to_integer(unsigned(andar_atual_in));
        destino_int := to_integer(unsigned(andar_destino_in));
        
        case estado_atual is
            
            when IDLE =>
                -- O elevador est� no andar de destino ou sem destino
                if atual_int /= destino_int then
                    -- H� um novo destino. Inicia o fechamento da porta.
                    proximo_estado <= FECHANDO_PORTA;
                    
                else 
                    -- N�o h� novo destino ou j� chegou. Fica em IDLE.
                    -- (Assumindo que em IDLE a porta pode estar aberta ou fechada)
                    proximo_estado <= IDLE;
                end if;
                
            when FECHANDO_PORTA =>
                start_close_out <= '1'; -- Sinaliza para a porta iniciar o fechamento
                
                if door_closed_in = '1' then
                    -- Porta fechou completamente (ap�s 2s, de acordo com porta.vhd)
                    proximo_estado <= MOVER;
                end if;

            when MOVER =>
                if atual_int /= destino_int then
                    motor_enable_out <= '1'; -- Liga o motor
                    
                    -- Define a dire��o do movimento
                    if direcao_req_in = '1' then -- Subir
                        move_up_out <= '1';
                    else                         -- Descer
                        move_down_out <= '1';
                    end if;
                    
                else
                    -- Chegou ao destino
                    proximo_estado <= CHEGOU_ANDAR;
                end if;
                
            when CHEGOU_ANDAR =>
                -- Para o motor (garantia, mesmo que j� estivesse parado)
                motor_enable_out <= '0';
                
                -- Limpa o bot�o que foi atendido (AQUI EST� A CHAVE)
                if botoes_pendentes_in(atual_int) = '1' then
                    -- Mant�m todos os outros bits, exceto o do andar atual
                    botoes_temp(atual_int) <= '0';
                end if;
                
                -- Ap�s limpar o pedido, a pr�xima a��o � abrir a porta
                proximo_estado <= ABRINDO_PORTA;
                
            when ABRINDO_PORTA =>
                -- Nenhuma a��o � necess�ria aqui. A porta permanece aberta (estado ABERTA em porta.vhd)
                
                -- Transi��o para o IDLE para aguardar novo destino ou fechamento de porta
                -- Para que o controlador n�o fique parado, volta para IDLE para verificar se h� um novo destino.
                proximo_estado <= IDLE; 
                
        end case;
    end process;
end architecture Behavioral;

