 --implementar depois :p